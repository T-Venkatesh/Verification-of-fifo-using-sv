`ifndef _bp_
`define _bp_

class basepkt;
bit wr;
bit rd;
rand bit [3:0]datain;
bit [3:0]dataout;
endclass
`endif    
